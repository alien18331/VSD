//================================================
// Auther:      Chang Wan-Yun (Claire)            
// Filename:    AXI.sv                            
// Description: Top module of AXI                  
// Version:     1.0 
//================================================
`include "AXI_define.svh"
`include "AR_Channel.sv"
`include "R_Channel.sv"
`include "AW_Channel.sv"
`include "W_Channel.sv"
`include "B_Channel.sv"


module AXI(

	input ACLK,
	input ARESETn,

	//SLAVE INTERFACE FOR MASTERS
	//WRITE ADDRESS
	input [`AXI_ID_BITS-1:0] AWID_M1,
	input [`AXI_ADDR_BITS-1:0] AWADDR_M1,
	input [`AXI_LEN_BITS-1:0] AWLEN_M1,
	input [`AXI_SIZE_BITS-1:0] AWSIZE_M1,
	input [1:0] AWBURST_M1,
	input AWVALID_M1,
	output AWREADY_M1,
	//WRITE DATA
	input [`AXI_DATA_BITS-1:0] WDATA_M1,
	input [`AXI_STRB_BITS-1:0] WSTRB_M1,
	input WLAST_M1,
	input WVALID_M1,
	output WREADY_M1,
	//WRITE RESPONSE
	output [`AXI_ID_BITS-1:0] BID_M1,
	output [3:0] BRESP_M1,
	output BVALID_M1,
	input BREADY_M1,
 
	//READ ADDRESS0
	input [`AXI_ID_BITS-1:0] ARID_M0,
	input [`AXI_ADDR_BITS-1:0] ARADDR_M0,
	input [`AXI_LEN_BITS-1:0] ARLEN_M0,
	input [`AXI_SIZE_BITS-1:0] ARSIZE_M0,
	input [1:0] ARBURST_M0,
	input ARVALID_M0,
	output ARREADY_M0,
	//READ DATA0
	output [`AXI_ID_BITS-1:0] RID_M0,
	output [`AXI_DATA_BITS-1:0] RDATA_M0,
	output [1:0] RRESP_M0,
	output RLAST_M0,
	output RVALID_M0,
	input RREADY_M0,
	//READ ADDRESS1
	input [`AXI_ID_BITS-1:0] ARID_M1,
	input [`AXI_ADDR_BITS-1:0] ARADDR_M1,
	input [`AXI_LEN_BITS-1:0] ARLEN_M1,
	input [`AXI_SIZE_BITS-1:0] ARSIZE_M1,
	input [1:0] ARBURST_M1,
	input ARVALID_M1,
	output ARREADY_M1,
	//READ DATA1
	output [`AXI_ID_BITS-1:0] RID_M1,
	output [`AXI_DATA_BITS-1:0] RDATA_M1,
	output [1:0] RRESP_M1,
	output RLAST_M1,
	output RVALID_M1,
	input RREADY_M1,

	//MASTER INTERFACE FOR SLAVES
	//WRITE ADDRESS0
	output [`AXI_IDS_BITS-1:0] AWID_S0,
	output [`AXI_ADDR_BITS-1:0] AWADDR_S0,
	output [`AXI_LEN_BITS-1:0] AWLEN_S0,
	output [`AXI_SIZE_BITS-1:0] AWSIZE_S0,
	output [1:0] AWBURST_S0,
	output AWVALID_S0,
	input AWREADY_S0,
	//WRITE DATA0
	output [`AXI_DATA_BITS-1:0] WDATA_S0,
	output [`AXI_STRB_BITS-1:0] WSTRB_S0,
	output WLAST_S0,
	output WVALID_S0,
	input WREADY_S0,
	//WRITE RESPONSE0
	input [`AXI_IDS_BITS-1:0] BID_S0,
	input [3:0] BRESP_S0,
	input BVALID_S0,
	output BREADY_S0,
	
	//WRITE ADDRESS1
	output [`AXI_IDS_BITS-1:0] AWID_S1,
	output [`AXI_ADDR_BITS-1:0] AWADDR_S1,
	output [`AXI_LEN_BITS-1:0] AWLEN_S1,
	output [`AXI_SIZE_BITS-1:0] AWSIZE_S1,
	output [1:0] AWBURST_S1,
	output AWVALID_S1,
	input AWREADY_S1,
	//WRITE DATA1
	output [`AXI_DATA_BITS-1:0] WDATA_S1,
	output [`AXI_STRB_BITS-1:0] WSTRB_S1,
	output WLAST_S1,
	output WVALID_S1,
	input WREADY_S1,
	//WRITE RESPONSE1
	input [`AXI_IDS_BITS-1:0] BID_S1,
	input [3:0] BRESP_S1,
	input BVALID_S1,
	output BREADY_S1,
	
	//READ ADDRESS0
	output [`AXI_IDS_BITS-1:0] ARID_S0,
	output [`AXI_ADDR_BITS-1:0] ARADDR_S0,
	output [`AXI_LEN_BITS-1:0] ARLEN_S0,
	output [`AXI_SIZE_BITS-1:0] ARSIZE_S0,
	output [1:0] ARBURST_S0,
	output ARVALID_S0,
	input ARREADY_S0,
	//READ DATA0
	input [`AXI_IDS_BITS-1:0] RID_S0,
	input [`AXI_DATA_BITS-1:0] RDATA_S0,
	input [1:0] RRESP_S0,
	input RLAST_S0,
	input RVALID_S0,
	output RREADY_S0,
	//READ ADDRESS1
	output [`AXI_IDS_BITS-1:0] ARID_S1,
	output [`AXI_ADDR_BITS-1:0] ARADDR_S1,
	output [`AXI_LEN_BITS-1:0] ARLEN_S1,
	output [`AXI_SIZE_BITS-1:0] ARSIZE_S1,
	output [1:0] ARBURST_S1,
	output ARVALID_S1,
	input ARREADY_S1,
	//READ DATA1
	input [`AXI_IDS_BITS-1:0] RID_S1,
	input [`AXI_DATA_BITS-1:0] RDATA_S1,
	input [1:0] RRESP_S1,
	input RLAST_S1,
	input RVALID_S1,
	output RREADY_S1
	
);
    //---------- you should put your design here ----------//
	
	logic R_done_M0;
	logic AR_R2S;
	logic [1:0] AW_W2S;
	logic [1:0] AW_W2S_0;
	// logic [1:0] W_done;
	
	AR_Channel AR(
		.clk(ACLK),
		.rst(~ARESETn),
		//READ ADDRESS0 - master0
		.ARID_M0(ARID_M0),
		.ARADDR_M0(ARADDR_M0),
		.ARLEN_M0(ARLEN_M0),
		.ARSIZE_M0(ARSIZE_M0),
		.ARBURST_M0(ARBURST_M0),
		.ARVALID_M0(ARVALID_M0),
		.ARREADY_M0(ARREADY_M0),
		//READ ADDRESS0 - master1
		.ARID_M1(ARID_M1),
		.ARADDR_M1(ARADDR_M1),
		.ARLEN_M1(ARLEN_M1),
		.ARSIZE_M1(ARSIZE_M1),
		.ARBURST_M1(ARBURST_M1),
		.ARVALID_M1(ARVALID_M1),
		.ARREADY_M1(ARREADY_M1),
		//READ ADDRESS0 - slave0
		.ARID_S0(ARID_S0),
		.ARADDR_S0(ARADDR_S0),
		.ARLEN_S0(ARLEN_S0),
		.ARSIZE_S0(ARSIZE_S0),
		.ARBURST_S0(ARBURST_S0),
		.ARVALID_S0(ARVALID_S0),
		.ARREADY_S0(ARREADY_S0),
		//READ ADDRESS0 - slave1
		.ARID_S1(ARID_S1),
		.ARADDR_S1(ARADDR_S1),
		.ARLEN_S1(ARLEN_S1),
		.ARSIZE_S1(ARSIZE_S1),
		.ARBURST_S1(ARBURST_S1),
		.ARVALID_S1(ARVALID_S1),
		.ARREADY_S1(ARREADY_S1),
		//From R_Channel
		.R_done_M0(R_done_M0),
		.R_done_M1(R_done_M1),
		.AR_R2S(AR_R2S)
	);
	
	R_Channel R(
		//READ DATA - slave0
		.RID_S0(RID_S0),
		.RDATA_S0(RDATA_S0),
		.RRESP_S0(RRESP_S0),
		.RLAST_S0(RLAST_S0),
		.RVALID_S0(RVALID_S0),
		.RREADY_S0(RREADY_S0),
		//READ DATA - slave1
		.RID_S1(RID_S1),
		.RDATA_S1(RDATA_S1),
		.RRESP_S1(RRESP_S1),
		.RLAST_S1(RLAST_S1),
		.RVALID_S1(RVALID_S1),
		.RREADY_S1(RREADY_S1),
		//READ DATA - master0
		.RID_M0(RID_M0),
		.RDATA_M0(RDATA_M0),
		.RRESP_M0(RRESP_M0),
		.RLAST_M0(RLAST_M0),
		.RVALID_M0(RVALID_M0),
		.RREADY_M0(RREADY_M0),
		//READ DATA - master1
		.RID_M1(RID_M1),
		.RDATA_M1(RDATA_M1),
		.RRESP_M1(RRESP_M1),
		.RLAST_M1(RLAST_M1),
		.RVALID_M1(RVALID_M1),
		.RREADY_M1(RREADY_M1),
		//AR_Channel
		.R_done_M0(R_done_M0),
		.R_done_M1(R_done_M1),
		.AR_R2S(AR_R2S)
	);
	
	AW_Channel AW(
		.clk(ACLK),
		.rst(~ARESETn),		
		//WRITE ADDRESS - master1
		.AWID_M1(AWID_M1),
		.AWADDR_M1(AWADDR_M1),
		.AWLEN_M1(AWLEN_M1),
		.AWSIZE_M1(AWSIZE_M1),
		.AWBURST_M1(AWBURST_M1),
		.AWVALID_M1(AWVALID_M1),
		.AWREADY_M1(AWREADY_M1),
		//WRITE ADDRESS - slave0
		.AWID_S0(AWID_S0),
		.AWADDR_S0(AWADDR_S0),
		.AWLEN_S0(AWLEN_S0),
		.AWSIZE_S0(AWSIZE_S0),
		.AWBURST_S0(AWBURST_S0),
		.AWVALID_S0(AWVALID_S0),
		.AWREADY_S0(AWREADY_S0),
		//WRITE ADDRESS - slave1
		.AWID_S1(AWID_S1),
		.AWADDR_S1(AWADDR_S1),
		.AWLEN_S1(AWLEN_S1),
		.AWSIZE_S1(AWSIZE_S1),
		.AWBURST_S1(AWBURST_S1),
		.AWVALID_S1(AWVALID_S1),
		.AWREADY_S1(AWREADY_S1),
		//W_Channel
		.AW_W2S(AW_W2S),
		.AW_W2S_0(AW_W2S_0),
		//B_Channel
		.B_done(B_done)
	);
	
	W_Channel W(
		.clk(ACLK),
		.rst(~ARESETn),
		//WRITE DATA - master1
		.WDATA_M1(WDATA_M1),
		.WSTRB_M1(WSTRB_M1),
		.WLAST_M1(WLAST_M1),
		.WVALID_M1(WVALID_M1),
		.WREADY_M1(WREADY_M1),
		//WRITE DATA - slave0
		.WDATA_S0(WDATA_S0),
		.WSTRB_S0(WSTRB_S0),
		.WLAST_S0(WLAST_S0),
		.WVALID_S0(WVALID_S0),
		.WREADY_S0(WREADY_S0),
		//WRITE DATA - slave1
		.WDATA_S1(WDATA_S1),
		.WSTRB_S1(WSTRB_S1),
		.WLAST_S1(WLAST_S1),
		.WVALID_S1(WVALID_S1),
		.WREADY_S1(WREADY_S1),
		//AW_Channel
		.AW_W2S(AW_W2S),
		.AW_W2S_0(AW_W2S_0),
		//B_Channel
		.B_done(B_done)	
	);
	
	B_Channel B(
		.clk(ACLK),
		.rst(~ARESETn),
		//WRITE RESPONSE - S0
		.BID_S0(BID_S0),
		.BRESP_S0(BRESP_S0),
		.BVALID_S0(BVALID_S0),
		.BREADY_S0(BREADY_S0),
		//WRITE RESPONSE - S1
		.BID_S1(BID_S1),
		.BRESP_S1(BRESP_S1),
		.BVALID_S1(BVALID_S1),
		.BREADY_S1(BREADY_S1),
		//WRITE RESPONSE - M0
		.BID_M0(),
		.BRESP_M0(),
		.BVALID_M0(),
		.BREADY_M0(1'b0),
		//WRITE RESPONSE - M1
		.BID_M1(BID_M1),
		.BRESP_M1(BRESP_M1),
		.BVALID_M1(BVALID_M1),
		.BREADY_M1(BREADY_M1),
		//B_Channel
		.B_done(B_done)
	);
	
	
	
endmodule
